

`define LANE_WIDTH 16
`define ADC_WIDTH 6
`define WAY_WIDTH 64
`define DES_OUT_WIDTH 4
`define DES_IN_WIDTH 2
`define PRLL_RANK 64
