

typedef struct packed {
  logic dpre;
  logic dpst;
  logic dcomp;
  logic dxp;
  logic dxn;
} ari_unit_t;

typedef struct packed {
  logic p1a;
  logic p1b;
  logic p2;
  logic p3o;
  logic p3a;
  logic p3b;
  logic p4p;
  logic p4m;
} flag_unit_t;
