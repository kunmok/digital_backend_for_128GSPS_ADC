

module scan_clkgen (
    RefClk,
    Reset,
    ClkEn,
    SClkP,
    SClkN
);

  //-----------------------------------------------------------------------------------
  //    System Inputs
  //-----------------------------------------------------------------------------------
  input wire RefClk;
  input wire Reset;
  input wire ClkEn;
  //-----------------------------------------------------------------------------------

  //-----------------------------------------------------------------------------------
  //    Outputs
  //-----------------------------------------------------------------------------------
  output wire SClkP;
  output wire SClkN;
  //-----------------------------------------------------------------------------------

  //-----------------------------------------------------------------------------------
  //    Signals
  //-----------------------------------------------------------------------------------
  reg [3:0] ShiftCountN;
  reg [3:0] ShiftCountP;
  //-----------------------------------------------------------------------------------

  //-----------------------------------------------------------------------------------
  //    Clock Generation
  //-----------------------------------------------------------------------------------
  assign SClkP = ShiftCountP[0];
  assign SClkN = ShiftCountN[0];
  //-----------------------------------------------------------------------------------

  //-----------------------------------------------------------------------------------
  //    Clock Generation
  //-----------------------------------------------------------------------------------
  always @(posedge RefClk or posedge Reset) begin
    if (Reset) ShiftCountP <= 4'b1000;
    else if (ClkEn) ShiftCountP <= {ShiftCountP[0], ShiftCountP[3:1]};
  end

  always @(posedge RefClk or posedge Reset) begin
    if (Reset) ShiftCountN <= 4'b0010;
    else if (ClkEn) ShiftCountN <= {ShiftCountN[0], ShiftCountN[3:1]};
  end
  //-----------------------------------------------------------------------------------

endmodule
