// updated LUT default table -> MSB is flipped to convert from unsigned binary to 2's complement format. 
`define LUT_DEFAULT_TABLE \
  { \
    6'b100000, \
    6'b100001, \
    6'b100010, \
    6'b100011, \
    6'b100100, \
    6'b100101, \
    6'b100110, \
    6'b100111, \
    6'b101100, \
    6'b101101, \
    6'b101110, \
    6'b101111, \
    6'b101000, \
    6'b101001, \
    6'b101010, \
    6'b101011, \
    6'b110000, \
    6'b110001, \
    6'b110010, \
    6'b110011, \
    6'b110100, \
    6'b110101, \
    6'b110110, \
    6'b110111, \
    6'b111100, \
    6'b111101, \
    6'b111110, \
    6'b111111, \
    6'b111000, \
    6'b111001, \
    6'b111010, \
    6'b111011, \
    6'b010000, \
    6'b010001, \
    6'b010010, \
    6'b010011, \
    6'b010100, \
    6'b010101, \
    6'b010110, \
    6'b010111, \
    6'b011100, \
    6'b011101, \
    6'b011110, \
    6'b011111, \
    6'b011000, \
    6'b011001, \
    6'b011010, \
    6'b011011, \
    6'b000000, \
    6'b000001, \
    6'b000010, \
    6'b000011, \
    6'b000100, \
    6'b000101, \
    6'b000110, \
    6'b000111, \
    6'b001100, \
    6'b001101, \
    6'b001110, \
    6'b001111, \
    6'b001000, \
    6'b001001, \
    6'b001010, \
    6'b001011 \
  }

// Lane physical-to-logical ordering (from bottom to top)
// 0 -> 8 -> 12 -> 4 -> 13 -> 5 -> 9 -> 1 -> 15 -> 7 -> 11 -> 3 -> 14 -> 6 -> 10 -> 2
`define LANE_PHYSICAL_ORDER '{0, 8, 12, 4, 13, 5, 9, 1, 15, 7, 11, 3, 14, 6, 10, 2}

`define DES_TO_LUT_PIPELINE_DEPTH 3
`define LUT_PIPELINE_DEPTH 1
`define REORDER_PIPELINE_DEPTH 4
