//==============================================================================
// Author: Sunjin Choi
// Description: 
// Signals:
// Note: 
// Variable naming conventions:
//    signals => snake_case
//    Parameters (aliasing signal values) => SNAKE_CASE with all caps
//    Parameters (not aliasing signal values) => CamelCase
//==============================================================================

// verilog_format: off
`timescale 1ns/1ps
`default_nettype none
// verilog_format: on

module pipeline_ff #(

) (

    // input signals

    // output signals

);

  // ----------------------------------------------------------------------
  // Parameters
  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------
  // Local Parameters
  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------
  // Inputs / Outputs
  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------
  // Signals
  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------
  // Assigns
  // ----------------------------------------------------------------------

  // ----------------------------------------------------------------------


endmodule

`default_nettype wire



