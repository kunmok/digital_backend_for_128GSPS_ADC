

/*`define NUM_BANKS 4
 *`define BANK_DEPTH 32*/

`define NUM_BANKS 8
`define BANK_DEPTH 16
`define MEM_WIDTH 384
`define FRAME_LENGTH 64
