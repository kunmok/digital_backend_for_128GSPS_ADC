
`timescale 1ns/1ps

// A bit-error-rate backend that supports counting the number of 1s (used for statistical eye)
// and for counting the number of bit-errors (used for BER eye)

module ber(
        clk,
        reset,

        mode,
        enable,
        
        in_test,
        in_correct,
        
        ber_count
    );

    //-----------------------------------------------------------------------------------
    //  Parameters
    //-----------------------------------------------------------------------------------
    parameter InWidth =             4;
    parameter CountWidth =          41;
    //-----------------------------------------------------------------------------------
    
    //-----------------------------------------------------------------------------------
    //  Constants
    //-----------------------------------------------------------------------------------
    localparam MWidth =             `log2(InWidth + 1);
    
    localparam Mode_Ones =          1'b0;
    localparam Mode_BER =           1'b1;
    //-----------------------------------------------------------------------------------

    //-----------------------------------------------------------------------------------
    //  I/O
    //-----------------------------------------------------------------------------------
    input wire                      clk;
    input wire                      reset;

    input wire                      mode;
    input wire                      enable;
    
    input wire  [InWidth-1:0]       in_test;
    input wire  [InWidth-1:0]       in_correct;
    
    output wire [CountWidth-1:0]    ber_count;
    //-----------------------------------------------------------------------------------

    //-----------------------------------------------------------------------------------
    //  Variables
    //-----------------------------------------------------------------------------------
    integer i;
    //-----------------------------------------------------------------------------------

    //-----------------------------------------------------------------------------------
    //  Signals
    //-----------------------------------------------------------------------------------
    reg         [MWidth-1:0]    mid_ctr, next_mid_ctr;
    wire        [InWidth-1:0]   errors;
    //-----------------------------------------------------------------------------------
            
    //-----------------------------------------------------------------------------------
    //  Assigns
    //-----------------------------------------------------------------------------------
    assign errors =             (mode == Mode_BER) ? in_test ^ in_correct : in_test;
    //-----------------------------------------------------------------------------------

    //-----------------------------------------------------------------------------------
    //  Intermediate Errors Counter
    //-----------------------------------------------------------------------------------
    // Sum up all errors in intermediate step
    always @(*) begin
        next_mid_ctr = {MWidth{1'b0}};
        if (enable) begin
            for (i = 0; i < InWidth; i = i + 1)
                next_mid_ctr = next_mid_ctr + errors[i];                
        end
    end

    always @ (posedge clk or posedge reset) begin
        if (reset) mid_ctr <= {MWidth{1'b0}};
        else mid_ctr <= next_mid_ctr;
    end
    //-----------------------------------------------------------------------------------
    
    //-----------------------------------------------------------------------------------
    //  Bit Errors Counter
    //-----------------------------------------------------------------------------------
    hybrid_counter  #   (   .Width      (CountWidth),
                            .SyncWidth  (MWidth))
            bit_counter (   .clk        (clk),
                            .reset      (reset),
                            .step       (mid_ctr),
                            .count      (ber_count));
    //-----------------------------------------------------------------------------------

    

endmodule

